//Release 2016.10.08
//File         : Processor_Pkg.sv
//Creator(s)   : Yang, Yu-Xiang (M10412034@yuntech.edu.tw)
//
//Description  : About Processor Port information  
//version : 1.0
//
package Processor_Pkg;



endpackage
